module fa(
input a , b, cin,
output co ,s 
);

ha ha1(a,b,co1,s1);
ha ha2(s1,cin,co2,s);
or or1(co,co1,co2);

endmodule